/*******************************************************
 * Copyright (C) 2022 German Iangalin, Bauman Moscow State Technical University,
 * Faculty of Rocket and Space Engineering.
 * All Rights Reserved.
 *
 * This file is part of  miriscv core.
 *
 *
 *******************************************************/

package  miriscv_cu_pkg;

  parameter NO_BYPASS = 2'd0;
  parameter BYPASS_E  = 2'd1;
  parameter BYPASS_M  = 2'd2;
  parameter BYPASS_W  = 2'd3;


endpackage :  miriscv_cu_pkg
